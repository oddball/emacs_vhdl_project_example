architecture rtl of block_bb is

begin




  

end architecture rtl;
