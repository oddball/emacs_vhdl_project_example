library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.projectname_components.all;

entity block_b is
  port (
    rstn : in std_ulogic;
    clk  : in std_ulogic);
end entity block_b;
