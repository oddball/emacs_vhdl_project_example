architecture rtl of block_aa is

begin

  

end architecture rtl;
